magic
tech sky130A
magscale 1 2
timestamp 1725542515
<< pwell >>
rect 3930 -190 4000 50
rect 4120 -190 4190 50
rect 4320 -190 4390 50
rect 4510 -190 4580 50
rect 4700 -190 4770 50
<< locali >>
rect 3930 3060 4770 3070
<< viali >>
rect 3230 3070 3390 3110
rect 3930 3070 4770 3110
rect 3220 -380 3400 -330
rect 3950 -370 4780 -330
<< metal1 >>
rect 2800 3320 4920 3480
rect 2800 3160 3940 3320
rect 4780 3160 4920 3320
rect 2800 3110 4920 3160
rect 2800 3070 3230 3110
rect 3390 3070 3930 3110
rect 4770 3070 4920 3110
rect 2800 3060 4920 3070
rect 3060 2920 3200 3060
rect 3280 2960 3360 3000
rect 3640 2960 4760 3000
rect 3640 2920 3800 2960
rect 3060 1120 3280 2920
rect 3340 1120 3800 2920
rect 3940 2920 4000 2930
rect 3940 2400 4000 2410
rect 4130 2920 4190 2930
rect 4130 2400 4190 2410
rect 4320 2920 4380 2930
rect 4320 2400 4380 2410
rect 4510 2920 4570 2930
rect 4510 2400 4570 2410
rect 4710 2920 4770 2930
rect 4710 2400 4770 2410
rect 4030 1640 4100 1650
rect 4030 1130 4100 1140
rect 4220 1640 4290 1650
rect 4220 1130 4290 1140
rect 4420 1640 4490 1650
rect 4420 1130 4490 1140
rect 4610 1640 4680 1650
rect 4610 1130 4680 1140
rect 2790 800 3020 870
rect 3280 800 3340 1080
rect 2790 660 3340 800
rect 2790 600 3020 660
rect 3280 440 3340 660
rect 3520 800 3800 1120
rect 3980 800 4760 1060
rect 4980 850 5210 870
rect 3520 660 4760 800
rect 4830 840 5210 850
rect 4830 690 4840 840
rect 4960 690 5210 840
rect 4830 670 5210 690
rect 3520 400 3800 660
rect 3980 460 4760 660
rect 4980 600 5210 670
rect 3040 -180 3280 400
rect 3340 -180 3800 400
rect 4030 370 4100 380
rect 4030 140 4100 150
rect 4220 370 4290 380
rect 4220 140 4290 150
rect 4420 370 4490 380
rect 4420 140 4490 150
rect 4610 370 4680 380
rect 4610 140 4680 150
rect 3040 -320 3200 -180
rect 3620 -220 3800 -180
rect 3930 40 4000 50
rect 3930 -190 4000 -180
rect 4120 40 4190 50
rect 4120 -190 4190 -180
rect 4320 40 4390 50
rect 4320 -190 4390 -180
rect 4510 40 4580 50
rect 4510 -190 4580 -180
rect 4700 40 4770 50
rect 4700 -190 4770 -180
rect 3280 -260 3360 -220
rect 3620 -260 4680 -220
rect 2800 -330 4920 -320
rect 2800 -380 3220 -330
rect 3400 -370 3950 -330
rect 4780 -370 4920 -330
rect 3400 -380 4920 -370
rect 2800 -390 4920 -380
rect 2800 -530 3940 -390
rect 4780 -530 4920 -390
rect 2800 -640 4920 -530
<< via1 >>
rect 3940 3160 4780 3320
rect 3940 2410 4000 2920
rect 4130 2410 4190 2920
rect 4320 2410 4380 2920
rect 4510 2410 4570 2920
rect 4710 2410 4770 2920
rect 4030 1140 4100 1640
rect 4220 1140 4290 1640
rect 4420 1140 4490 1640
rect 4610 1140 4680 1640
rect 4840 690 4960 840
rect 4030 150 4100 370
rect 4220 150 4290 370
rect 4420 150 4490 370
rect 4610 150 4680 370
rect 3930 -180 4000 40
rect 4120 -180 4190 40
rect 4320 -180 4390 40
rect 4510 -180 4580 40
rect 4700 -180 4770 40
rect 3940 -530 4780 -390
<< metal2 >>
rect 3920 3320 4800 3340
rect 3920 3160 3940 3320
rect 4780 3160 4800 3320
rect 3920 2920 4800 3160
rect 3920 2410 3940 2920
rect 4000 2410 4130 2920
rect 4190 2410 4320 2920
rect 4380 2410 4510 2920
rect 4570 2410 4710 2920
rect 4770 2410 4800 2920
rect 3920 2360 4800 2410
rect 3920 1640 4800 1680
rect 3920 1140 4030 1640
rect 4100 1140 4220 1640
rect 4290 1140 4420 1640
rect 4490 1140 4610 1640
rect 4680 1140 4800 1640
rect 3920 890 4800 1140
rect 3920 840 4970 890
rect 3920 690 4840 840
rect 4960 690 4970 840
rect 3920 630 4970 690
rect 3920 370 4800 630
rect 3920 150 4030 370
rect 4100 150 4220 370
rect 4290 150 4420 370
rect 4490 150 4610 370
rect 4680 150 4800 370
rect 3920 130 4800 150
rect 3920 40 4800 60
rect 3920 -180 3930 40
rect 4000 -180 4120 40
rect 4190 -180 4320 40
rect 4390 -180 4510 40
rect 4580 -180 4700 40
rect 4770 -180 4800 40
rect 3920 -390 4800 -180
rect 3920 -530 3940 -390
rect 4780 -530 4800 -390
rect 3920 -550 4800 -530
use sky130_fd_pr__pfet_01v8_XGSFBL  XM9
timestamp 1725540246
transform 1 0 3311 0 1 2019
box -211 -1119 211 1119
use sky130_fd_pr__nfet_01v8_J2SMEF  XM10
timestamp 1725540246
transform 1 0 3311 0 1 110
box -211 -510 211 510
use sky130_fd_pr__pfet_01v8_UG67RG  XM11
timestamp 1725540246
transform 1 0 4351 0 1 2019
box -551 -1119 551 1119
use sky130_fd_pr__nfet_01v8_F5PS5H  XM12
timestamp 1725540246
transform 1 0 4351 0 1 110
box -551 -510 551 510
<< labels >>
flabel metal1 2800 600 3000 800 0 FreeSans 256 0 0 0 in
port 2 nsew
flabel metal1 5000 600 5200 800 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 2800 3280 3000 3480 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 2800 -640 3000 -440 0 FreeSans 256 0 0 0 VSS
port 1 nsew
<< end >>
