magic
tech sky130A
timestamp 1725622005
<< metal2 >>
rect 756 2492 784 2520
rect 7728 2492 7756 2520
rect 756 2464 840 2492
rect 4312 2464 4368 2492
rect 7728 2464 7812 2492
rect 756 2436 896 2464
rect 4312 2436 4424 2464
rect 7728 2436 7840 2464
rect 756 2408 952 2436
rect 4312 2408 4480 2436
rect 7728 2408 7924 2436
rect 756 2380 1008 2408
rect 4312 2380 4536 2408
rect 7728 2380 7980 2408
rect 756 2352 1064 2380
rect 4312 2352 4592 2380
rect 7728 2352 8008 2380
rect 756 2324 1120 2352
rect 4312 2324 4648 2352
rect 7728 2324 8092 2352
rect 756 1680 868 2324
rect 924 2296 1176 2324
rect 980 2268 1232 2296
rect 1036 2240 1288 2268
rect 1092 2212 1344 2240
rect 1148 2184 1400 2212
rect 1204 2156 1456 2184
rect 1260 2128 1512 2156
rect 1316 2100 1568 2128
rect 1372 2072 1624 2100
rect 1428 2044 1680 2072
rect 1484 2016 1736 2044
rect 1540 1988 1792 2016
rect 1596 1960 1848 1988
rect 1652 1932 1904 1960
rect 1708 1904 1960 1932
rect 1764 1876 2016 1904
rect 1820 1848 2072 1876
rect 1876 1820 2128 1848
rect 1932 1792 2184 1820
rect 2436 1792 2576 1820
rect 1988 1764 2240 1792
rect 2380 1764 2632 1792
rect 2044 1736 2296 1764
rect 2352 1736 2660 1764
rect 2100 1708 2436 1736
rect 2576 1708 2688 1736
rect 2156 1680 2408 1708
rect 2604 1680 2688 1708
rect 4312 1680 4424 2324
rect 4452 2296 4704 2324
rect 4508 2268 4760 2296
rect 4564 2240 4816 2268
rect 4620 2212 4872 2240
rect 4676 2184 4928 2212
rect 4732 2156 4984 2184
rect 4788 2128 5040 2156
rect 4844 2100 5096 2128
rect 4900 2072 5152 2100
rect 4956 2044 5208 2072
rect 5040 2016 5264 2044
rect 5068 1988 5320 2016
rect 5124 1960 5376 1988
rect 5208 1932 5432 1960
rect 5236 1904 5488 1932
rect 5292 1876 5544 1904
rect 5376 1848 5600 1876
rect 5404 1820 5684 1848
rect 5460 1792 5712 1820
rect 5964 1792 6132 1820
rect 5544 1764 5768 1792
rect 5936 1764 6188 1792
rect 5572 1736 5852 1764
rect 5908 1736 6216 1764
rect 5628 1708 5964 1736
rect 6132 1708 6216 1736
rect 5712 1680 5936 1708
rect 0 1596 868 1680
rect 2212 1652 2380 1680
rect 2268 1624 2380 1652
rect 2240 1596 2380 1624
rect 2632 1596 4424 1680
rect 5740 1652 5936 1680
rect 6160 1680 6244 1708
rect 7728 1680 7840 2324
rect 7896 2296 8148 2324
rect 7952 2268 8176 2296
rect 8008 2240 8260 2268
rect 8064 2212 8316 2240
rect 8120 2184 8344 2212
rect 8176 2156 8428 2184
rect 8232 2128 8484 2156
rect 8288 2100 8540 2128
rect 8344 2072 8596 2100
rect 8400 2044 8652 2072
rect 8456 2016 8708 2044
rect 8512 1988 8764 2016
rect 8568 1960 8820 1988
rect 8624 1932 8876 1960
rect 8680 1904 8932 1932
rect 8736 1876 8988 1904
rect 8792 1848 9044 1876
rect 8848 1820 9100 1848
rect 8904 1792 9156 1820
rect 9408 1792 9548 1820
rect 8960 1764 9212 1792
rect 9352 1764 9604 1792
rect 9016 1736 9268 1764
rect 9324 1736 9632 1764
rect 10836 1736 10864 1764
rect 9072 1708 9380 1736
rect 9548 1708 9632 1736
rect 10332 1708 10472 1736
rect 10836 1708 10948 1736
rect 9128 1680 9380 1708
rect 9576 1680 9660 1708
rect 10304 1680 10500 1708
rect 10836 1680 11088 1708
rect 6160 1652 7840 1680
rect 9184 1652 9352 1680
rect 5796 1596 5936 1652
rect 6188 1624 7840 1652
rect 9240 1624 9352 1652
rect 0 84 84 1596
rect 756 952 868 1596
rect 2184 1568 2408 1596
rect 2632 1568 2688 1596
rect 2128 1540 2408 1568
rect 2604 1540 2688 1568
rect 2072 1512 2436 1540
rect 2576 1512 2660 1540
rect 2016 1484 2268 1512
rect 2352 1484 2660 1512
rect 1960 1456 2212 1484
rect 2408 1456 2632 1484
rect 1904 1428 2156 1456
rect 2464 1428 2548 1456
rect 1848 1400 2100 1428
rect 1792 1372 2044 1400
rect 1736 1344 1988 1372
rect 1680 1316 1932 1344
rect 1624 1288 1876 1316
rect 1568 1260 1820 1288
rect 1512 1232 1764 1260
rect 1456 1204 1708 1232
rect 1400 1176 1652 1204
rect 1344 1148 1596 1176
rect 1288 1120 1540 1148
rect 1232 1092 1484 1120
rect 1176 1064 1428 1092
rect 1120 1036 1372 1064
rect 1064 1008 1316 1036
rect 1008 980 1260 1008
rect 952 952 1204 980
rect 4312 952 4424 1596
rect 5740 1568 5936 1596
rect 6160 1596 7840 1624
rect 9212 1596 9352 1624
rect 9604 1596 11200 1680
rect 5684 1540 5964 1568
rect 6160 1540 6244 1596
rect 5628 1512 5992 1540
rect 6104 1512 6216 1540
rect 5572 1484 5824 1512
rect 5908 1484 6188 1512
rect 5516 1456 5768 1484
rect 5936 1456 6160 1484
rect 5460 1428 5712 1456
rect 5992 1428 6104 1456
rect 5404 1400 5656 1428
rect 5348 1372 5600 1400
rect 5292 1344 5544 1372
rect 5236 1316 5488 1344
rect 5180 1288 5432 1316
rect 5124 1260 5376 1288
rect 5068 1232 5320 1260
rect 5012 1204 5264 1232
rect 4956 1176 5208 1204
rect 4900 1148 5152 1176
rect 4844 1120 5096 1148
rect 4788 1092 5040 1120
rect 4732 1064 4984 1092
rect 4676 1036 4900 1064
rect 4620 1008 4872 1036
rect 4564 980 4816 1008
rect 4508 952 4732 980
rect 7728 952 7840 1596
rect 9156 1568 9352 1596
rect 9100 1540 9380 1568
rect 9576 1540 9660 1596
rect 10276 1568 10500 1596
rect 10836 1568 11172 1596
rect 10304 1540 10472 1568
rect 10836 1540 11032 1568
rect 9044 1512 9408 1540
rect 9548 1512 9632 1540
rect 10332 1512 10444 1540
rect 10836 1512 10920 1540
rect 8988 1484 9240 1512
rect 9324 1484 9632 1512
rect 8932 1456 9184 1484
rect 9352 1456 9576 1484
rect 8876 1428 9128 1456
rect 9436 1428 9520 1456
rect 8820 1400 9072 1428
rect 8764 1372 9016 1400
rect 8708 1344 8960 1372
rect 8652 1316 8904 1344
rect 8596 1288 8848 1316
rect 8540 1260 8792 1288
rect 8484 1232 8736 1260
rect 8428 1204 8680 1232
rect 8372 1176 8624 1204
rect 8316 1148 8568 1176
rect 8260 1120 8512 1148
rect 8204 1092 8456 1120
rect 8148 1064 8400 1092
rect 8092 1036 8344 1064
rect 8036 1008 8288 1036
rect 7980 980 8232 1008
rect 7924 952 8176 980
rect 756 924 1148 952
rect 4312 924 4704 952
rect 7728 924 8120 952
rect 756 896 1092 924
rect 4312 896 4648 924
rect 7728 896 8064 924
rect 756 868 1036 896
rect 4312 868 4564 896
rect 7728 868 8008 896
rect 756 840 980 868
rect 4312 840 4536 868
rect 7728 840 7952 868
rect 756 812 924 840
rect 4312 812 4480 840
rect 7728 812 7896 840
rect 756 784 868 812
rect 4312 784 4424 812
rect 7728 784 7840 812
rect 756 756 812 784
rect 4312 756 4368 784
rect 7728 756 7784 784
rect 10360 84 10444 1512
rect 0 0 10444 84
<< end >>
