magic
tech sky130A
magscale 1 2
timestamp 1725540246
<< error_p >>
rect -29 981 29 987
rect -29 947 -17 981
rect -29 941 29 947
rect -29 -947 29 -941
rect -29 -981 -17 -947
rect -29 -987 29 -981
<< nwell >>
rect -211 -1119 211 1119
<< pmos >>
rect -15 -900 15 900
<< pdiff >>
rect -73 888 -15 900
rect -73 -888 -61 888
rect -27 -888 -15 888
rect -73 -900 -15 -888
rect 15 888 73 900
rect 15 -888 27 888
rect 61 -888 73 888
rect 15 -900 73 -888
<< pdiffc >>
rect -61 -888 -27 888
rect 27 -888 61 888
<< nsubdiff >>
rect -175 1049 -79 1083
rect 79 1049 175 1083
rect -175 987 -141 1049
rect 141 987 175 1049
rect -175 -1049 -141 -987
rect 141 -1049 175 -987
rect -175 -1083 -79 -1049
rect 79 -1083 175 -1049
<< nsubdiffcont >>
rect -79 1049 79 1083
rect -175 -987 -141 987
rect 141 -987 175 987
rect -79 -1083 79 -1049
<< poly >>
rect -33 981 33 997
rect -33 947 -17 981
rect 17 947 33 981
rect -33 931 33 947
rect -15 900 15 931
rect -15 -931 15 -900
rect -33 -947 33 -931
rect -33 -981 -17 -947
rect 17 -981 33 -947
rect -33 -997 33 -981
<< polycont >>
rect -17 947 17 981
rect -17 -981 17 -947
<< locali >>
rect -175 1049 -79 1083
rect 79 1049 175 1083
rect -175 987 -141 1049
rect 141 987 175 1049
rect -33 947 -17 981
rect 17 947 33 981
rect -61 888 -27 904
rect -61 -904 -27 -888
rect 27 888 61 904
rect 27 -904 61 -888
rect -33 -981 -17 -947
rect 17 -981 33 -947
rect -175 -1049 -141 -987
rect 141 -1049 175 -987
rect -175 -1083 -79 -1049
rect 79 -1083 175 -1049
<< viali >>
rect -17 947 17 981
rect -61 -888 -27 888
rect 27 -888 61 888
rect -17 -981 17 -947
<< metal1 >>
rect -29 981 29 987
rect -29 947 -17 981
rect 17 947 29 981
rect -29 941 29 947
rect -67 888 -21 900
rect -67 -888 -61 888
rect -27 -888 -21 888
rect -67 -900 -21 -888
rect 21 888 67 900
rect 21 -888 27 888
rect 61 -888 67 888
rect 21 -900 67 -888
rect -29 -947 29 -941
rect -29 -981 -17 -947
rect 17 -981 29 -947
rect -29 -987 29 -981
<< properties >>
string FIXED_BBOX -158 -1066 158 1066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
