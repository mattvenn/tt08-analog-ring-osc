magic
tech sky130A
magscale 1 2
timestamp 1725561279
<< metal1 >>
rect 27794 7440 27800 7840
rect 28200 7440 28700 7840
rect 29920 7180 30760 7540
rect 29900 6780 30260 6800
rect 27760 6500 29480 6780
rect 29900 6500 29940 6780
rect 30220 6500 30260 6780
rect 27760 3340 28040 6500
rect 29900 6480 30260 6500
rect 28400 5680 28800 5920
rect 28394 5280 28400 5680
rect 28800 5280 28806 5680
rect 30400 5560 30760 7180
rect 27760 3060 28640 3340
rect 27874 1920 27880 2320
rect 28280 2280 28520 2320
rect 28280 1920 28540 2280
rect 28300 1800 28540 1920
rect 30610 1205 30820 3305
rect 30295 1090 30820 1205
rect 30295 995 30362 1090
rect 30356 910 30362 995
rect 30542 995 30820 1090
rect 30542 910 30548 995
<< via1 >>
rect 27800 7440 28200 7840
rect 29940 6500 30220 6780
rect 28400 5280 28800 5680
rect 27880 1920 28280 2320
rect 30362 910 30542 1090
<< metal2 >>
rect 30400 8740 30680 8749
rect 27800 7840 28200 7846
rect 27796 7440 27800 7495
rect 28200 7440 28204 7495
rect 27796 7105 27805 7440
rect 28195 7105 28204 7440
rect 27800 7100 28200 7105
rect 29900 6780 30260 6800
rect 30400 6780 30680 8460
rect 29900 6500 29940 6780
rect 30220 6500 30680 6780
rect 29900 6480 30260 6500
rect 28400 5680 28800 5686
rect 28400 5055 28800 5280
rect 28396 4665 28405 5055
rect 28795 4665 28804 5055
rect 28400 4660 28800 4665
rect 27880 2575 28280 2580
rect 27876 2320 27885 2575
rect 28275 2320 28284 2575
rect 27876 2185 27880 2320
rect 28280 2185 28284 2320
rect 27880 1914 28280 1920
rect 30362 1090 30542 1096
rect 30362 885 30542 910
rect 30358 715 30367 885
rect 30537 715 30546 885
rect 30362 710 30542 715
<< via2 >>
rect 30400 8460 30680 8740
rect 27805 7440 28195 7495
rect 27805 7105 28195 7440
rect 28405 4665 28795 5055
rect 27885 2320 28275 2575
rect 27885 2185 28275 2320
rect 30367 715 30537 885
<< metal3 >>
rect 30400 10040 30680 10046
rect 30400 8745 30680 9760
rect 30395 8740 30685 8745
rect 30395 8460 30400 8740
rect 30680 8460 30685 8740
rect 30395 8455 30685 8460
rect 27800 7495 28200 7500
rect 27800 7139 27805 7495
rect 28195 7139 28200 7495
rect 27795 6741 27801 7139
rect 28199 6741 28205 7139
rect 27800 6740 28200 6741
rect 28400 5055 28800 5060
rect 28400 4700 28405 5055
rect 200 4680 28405 4700
rect 200 4320 220 4680
rect 580 4665 28405 4680
rect 28795 4700 28800 5055
rect 28795 4665 30500 4700
rect 580 4320 30500 4665
rect 200 4300 30500 4320
rect 27880 2819 28280 2820
rect 27875 2421 27881 2819
rect 28279 2421 28285 2819
rect 27880 2185 27885 2421
rect 28275 2185 28280 2421
rect 27880 2180 28280 2185
rect 30362 885 30542 890
rect 30362 715 30367 885
rect 30537 715 30542 885
rect 30362 589 30542 715
rect 30357 411 30363 589
rect 30541 411 30547 589
rect 30362 410 30542 411
<< via3 >>
rect 30400 9760 30680 10040
rect 27801 7105 27805 7139
rect 27805 7105 28195 7139
rect 28195 7105 28199 7139
rect 27801 6741 28199 7105
rect 220 4320 580 4680
rect 27881 2575 28279 2819
rect 27881 2421 27885 2575
rect 27885 2421 28275 2575
rect 28275 2421 28279 2575
rect 30363 411 30541 589
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 200 4680 600 44152
rect 200 4320 220 4680
rect 580 4320 600 4680
rect 200 1000 600 4320
rect 800 5500 1200 44152
rect 27662 43370 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 30400 43370 30680 43400
rect 27662 43310 30680 43370
rect 30400 10041 30680 43310
rect 30399 10040 30681 10041
rect 30399 9760 30400 10040
rect 30680 9760 30681 10040
rect 30399 9759 30681 9760
rect 27800 7139 28200 7140
rect 27800 6741 27801 7139
rect 28199 6741 28200 7139
rect 27800 5500 28200 6741
rect 800 5100 30600 5500
rect 800 1000 1200 5100
rect 27880 2819 28280 5100
rect 27880 2421 27881 2819
rect 28279 2421 28280 2819
rect 27880 2420 28280 2421
rect 30362 589 30542 590
rect 30362 411 30363 589
rect 30541 411 30542 589
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 411
use driver  driver_0 ~/work/asic-workshop/shuttle-tt08/tt08-analog-ring-osc/mag
timestamp 1725547227
transform 1 0 25610 0 1 2440
box 2790 -640 5210 3480
use ring  ring_0
timestamp 1725561279
transform 0 1 29640 -1 0 11140
box -220 -1240 4640 640
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
