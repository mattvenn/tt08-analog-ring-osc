magic
tech sky130A
timestamp 1725621121
<< metal2 >>
rect 1260 4144 1288 4172
rect 7112 4144 7140 4172
rect 12796 4144 12824 4172
rect 1260 4116 1344 4144
rect 7112 4116 7196 4144
rect 12768 4116 12880 4144
rect 1260 4088 1400 4116
rect 7112 4088 7252 4116
rect 12768 4088 12936 4116
rect 18200 4088 18228 4116
rect 1260 4060 1456 4088
rect 7112 4060 7308 4088
rect 12768 4060 12992 4088
rect 18060 4060 18368 4088
rect 1260 4032 1512 4060
rect 7112 4032 7364 4060
rect 12768 4032 13048 4060
rect 18004 4032 18200 4060
rect 18228 4032 18424 4060
rect 1260 4004 1568 4032
rect 7112 4004 7420 4032
rect 12768 4004 13076 4032
rect 17976 4004 18088 4032
rect 18340 4004 18452 4032
rect 1260 3976 1624 4004
rect 7112 3976 7476 4004
rect 12768 3976 13160 4004
rect 17920 3976 18032 4004
rect 18368 3976 18480 4004
rect 1260 3948 1680 3976
rect 7112 3948 7532 3976
rect 12768 3948 13216 3976
rect 17892 3948 18004 3976
rect 18396 3948 18480 3976
rect 1260 3920 1736 3948
rect 7112 3920 7588 3948
rect 12768 3920 13244 3948
rect 17864 3920 17976 3948
rect 1260 3892 1792 3920
rect 7112 3892 7644 3920
rect 12768 3892 13328 3920
rect 17864 3892 17948 3920
rect 1260 3864 1848 3892
rect 7112 3864 7700 3892
rect 12768 3864 13384 3892
rect 17836 3864 17948 3892
rect 18396 3864 18508 3948
rect 1260 3836 1904 3864
rect 7112 3836 7756 3864
rect 12768 3836 13412 3864
rect 1260 2772 1456 3836
rect 1512 3808 1960 3836
rect 1568 3780 2016 3808
rect 1624 3752 2072 3780
rect 1680 3724 2128 3752
rect 1736 3696 2184 3724
rect 1792 3668 2240 3696
rect 1848 3640 2296 3668
rect 1904 3612 2352 3640
rect 1960 3584 2408 3612
rect 2016 3556 2464 3584
rect 2072 3528 2520 3556
rect 2128 3500 2576 3528
rect 2184 3472 2632 3500
rect 2240 3444 2688 3472
rect 2296 3416 2744 3444
rect 2352 3388 2800 3416
rect 2408 3360 2856 3388
rect 2464 3332 2912 3360
rect 2520 3304 2968 3332
rect 2576 3276 3024 3304
rect 2632 3248 3080 3276
rect 2688 3220 3136 3248
rect 2744 3192 3192 3220
rect 2800 3164 3248 3192
rect 2856 3136 3304 3164
rect 2912 3108 3360 3136
rect 2968 3080 3416 3108
rect 3024 3052 3472 3080
rect 3080 3024 3528 3052
rect 3136 2996 3584 3024
rect 4060 2996 4256 3024
rect 3192 2968 3640 2996
rect 3976 2968 4312 2996
rect 3248 2940 3696 2968
rect 3948 2940 4340 2968
rect 3304 2912 3752 2940
rect 3920 2912 4396 2940
rect 3360 2884 3808 2912
rect 3892 2884 4396 2912
rect 3416 2856 4060 2884
rect 4256 2856 4424 2884
rect 3472 2828 4004 2856
rect 4284 2828 4452 2856
rect 3528 2800 4004 2828
rect 3584 2772 3976 2800
rect 4312 2772 4452 2828
rect 7112 2772 7308 3836
rect 7364 3808 7812 3836
rect 7420 3780 7868 3808
rect 7476 3752 7924 3780
rect 7532 3724 7980 3752
rect 7588 3696 8036 3724
rect 7644 3668 8092 3696
rect 7700 3640 8148 3668
rect 7756 3612 8204 3640
rect 7812 3584 8260 3612
rect 7868 3556 8316 3584
rect 7924 3528 8372 3556
rect 7980 3500 8428 3528
rect 8036 3472 8484 3500
rect 8092 3444 8540 3472
rect 8148 3416 8596 3444
rect 8204 3388 8652 3416
rect 8260 3360 8708 3388
rect 8316 3332 8764 3360
rect 8372 3304 8820 3332
rect 8428 3276 8876 3304
rect 8484 3248 8932 3276
rect 8540 3220 8988 3248
rect 8596 3192 9044 3220
rect 8652 3164 9100 3192
rect 8736 3136 9156 3164
rect 8792 3108 9212 3136
rect 8848 3080 9268 3108
rect 8904 3052 9324 3080
rect 8960 3024 9380 3052
rect 9016 2996 9436 3024
rect 9912 2996 10108 3024
rect 9072 2968 9492 2996
rect 9856 2968 10164 2996
rect 9128 2940 9548 2968
rect 9800 2940 10220 2968
rect 9184 2912 9604 2940
rect 9772 2912 10248 2940
rect 9240 2884 9660 2912
rect 9744 2884 10276 2912
rect 9296 2856 9912 2884
rect 10108 2856 10304 2884
rect 9352 2828 9884 2856
rect 10136 2828 10304 2856
rect 9408 2800 9856 2828
rect 10164 2800 10332 2828
rect 9464 2772 9828 2800
rect 0 2632 1456 2772
rect 3640 2744 3976 2772
rect 3696 2716 3948 2744
rect 3752 2688 3948 2716
rect 3724 2660 3948 2688
rect 3668 2632 3948 2660
rect 4340 2632 7308 2772
rect 9520 2744 9828 2772
rect 10192 2772 10332 2800
rect 12768 2772 12992 3836
rect 13048 3808 13496 3836
rect 13104 3780 13552 3808
rect 17808 3780 17920 3864
rect 18396 3836 18536 3864
rect 18424 3808 18536 3836
rect 13160 3752 13608 3780
rect 13216 3724 13664 3752
rect 13272 3696 13720 3724
rect 13328 3668 13776 3696
rect 17780 3668 17892 3780
rect 13384 3640 13832 3668
rect 17752 3640 17892 3668
rect 18396 3752 18536 3808
rect 18396 3640 18508 3752
rect 13440 3612 13888 3640
rect 13496 3584 13944 3612
rect 13552 3556 14000 3584
rect 17752 3556 17864 3640
rect 18368 3612 18508 3640
rect 18368 3556 18480 3612
rect 13608 3528 14056 3556
rect 17752 3528 17892 3556
rect 13664 3500 14112 3528
rect 13720 3472 14168 3500
rect 13776 3444 14224 3472
rect 17780 3444 17892 3528
rect 18340 3500 18452 3556
rect 18312 3472 18424 3500
rect 18284 3444 18396 3472
rect 13832 3416 14280 3444
rect 17808 3416 17920 3444
rect 18256 3416 18368 3444
rect 13888 3388 14336 3416
rect 17836 3388 17948 3416
rect 18228 3388 18340 3416
rect 13944 3360 14392 3388
rect 17864 3360 18004 3388
rect 18172 3360 18284 3388
rect 14000 3332 14448 3360
rect 17892 3332 18256 3360
rect 14056 3304 14504 3332
rect 17976 3304 18172 3332
rect 14112 3276 14560 3304
rect 18088 3276 18172 3304
rect 14168 3248 14616 3276
rect 18088 3248 18228 3276
rect 14224 3220 14672 3248
rect 18116 3220 18424 3248
rect 14280 3192 14728 3220
rect 18144 3192 18424 3220
rect 14336 3164 14784 3192
rect 18200 3164 18424 3192
rect 14392 3136 14840 3164
rect 14448 3108 14896 3136
rect 14504 3080 14952 3108
rect 14560 3052 15008 3080
rect 14616 3024 15064 3052
rect 14672 2996 15120 3024
rect 15596 2996 15764 3024
rect 14728 2968 15176 2996
rect 15512 2968 15848 2996
rect 14784 2940 15232 2968
rect 15484 2940 15876 2968
rect 14840 2912 15288 2940
rect 15456 2912 15904 2940
rect 14896 2884 15344 2912
rect 15428 2884 15932 2912
rect 17920 2884 18004 2912
rect 14952 2856 15596 2884
rect 15764 2856 15960 2884
rect 17108 2856 17304 2884
rect 17920 2856 18116 2884
rect 15008 2828 15540 2856
rect 15820 2828 15988 2856
rect 17080 2828 17332 2856
rect 17920 2828 18228 2856
rect 15064 2800 15512 2828
rect 15120 2772 15512 2800
rect 15848 2772 15988 2828
rect 17052 2800 17360 2828
rect 17920 2800 18340 2828
rect 17024 2772 17388 2800
rect 17920 2772 18452 2800
rect 10192 2744 12992 2772
rect 15176 2744 15484 2772
rect 9576 2716 9828 2744
rect 9604 2688 9828 2716
rect 9576 2660 9828 2688
rect 10220 2660 12992 2744
rect 15232 2716 15484 2744
rect 15288 2688 15484 2716
rect 15260 2660 15484 2688
rect 9520 2632 9828 2660
rect 0 140 140 2632
rect 1260 1540 1456 2632
rect 3612 2604 3976 2632
rect 4340 2604 4480 2632
rect 3556 2576 3976 2604
rect 4312 2576 4452 2604
rect 3500 2548 4004 2576
rect 4284 2548 4452 2576
rect 3444 2520 4032 2548
rect 4256 2520 4424 2548
rect 3388 2492 3836 2520
rect 3892 2492 4116 2520
rect 4200 2492 4424 2520
rect 3332 2464 3780 2492
rect 3892 2464 4396 2492
rect 3276 2436 3724 2464
rect 3948 2436 4368 2464
rect 3220 2408 3668 2436
rect 3976 2408 4340 2436
rect 3164 2380 3612 2408
rect 4032 2380 4284 2408
rect 3108 2352 3556 2380
rect 3052 2324 3500 2352
rect 2996 2296 3444 2324
rect 2940 2268 3388 2296
rect 2884 2240 3332 2268
rect 2828 2212 3276 2240
rect 2772 2184 3220 2212
rect 2716 2156 3164 2184
rect 2660 2128 3108 2156
rect 2604 2100 3052 2128
rect 2548 2072 2996 2100
rect 2492 2044 2940 2072
rect 2436 2016 2884 2044
rect 2380 1988 2828 2016
rect 2324 1960 2772 1988
rect 2268 1932 2716 1960
rect 2212 1904 2660 1932
rect 2156 1876 2604 1904
rect 2100 1848 2548 1876
rect 2044 1820 2492 1848
rect 1988 1792 2436 1820
rect 1932 1764 2380 1792
rect 1876 1736 2324 1764
rect 1820 1708 2268 1736
rect 1764 1680 2212 1708
rect 1708 1652 2156 1680
rect 1652 1624 2100 1652
rect 1596 1596 2044 1624
rect 1540 1568 1988 1596
rect 1484 1540 1904 1568
rect 7112 1540 7308 2632
rect 9464 2604 9828 2632
rect 10192 2632 12992 2660
rect 15204 2632 15484 2660
rect 15876 2632 18536 2772
rect 9408 2576 9856 2604
rect 10192 2576 10332 2632
rect 9352 2548 9884 2576
rect 10164 2548 10304 2576
rect 9296 2520 9912 2548
rect 10136 2520 10304 2548
rect 9240 2492 9688 2520
rect 9744 2492 9968 2520
rect 10052 2492 10276 2520
rect 9184 2464 9632 2492
rect 9772 2464 10248 2492
rect 9128 2436 9576 2464
rect 9800 2436 10220 2464
rect 9072 2408 9520 2436
rect 9828 2408 10192 2436
rect 9016 2380 9464 2408
rect 9884 2380 10136 2408
rect 8960 2352 9408 2380
rect 8904 2324 9352 2352
rect 8848 2296 9296 2324
rect 8792 2268 9240 2296
rect 8736 2240 9184 2268
rect 8680 2212 9128 2240
rect 8624 2184 9072 2212
rect 8568 2156 9016 2184
rect 8512 2128 8960 2156
rect 8456 2100 8904 2128
rect 8400 2072 8848 2100
rect 8344 2044 8792 2072
rect 8288 2016 8736 2044
rect 8232 1988 8680 2016
rect 8176 1960 8624 1988
rect 8120 1932 8568 1960
rect 8064 1904 8512 1932
rect 8008 1876 8456 1904
rect 7952 1848 8400 1876
rect 7896 1820 8344 1848
rect 7840 1792 8288 1820
rect 7784 1764 8232 1792
rect 7728 1736 8176 1764
rect 7672 1708 8120 1736
rect 7616 1680 8064 1708
rect 7560 1652 8008 1680
rect 7504 1624 7952 1652
rect 7448 1596 7896 1624
rect 7392 1568 7840 1596
rect 12768 1568 12992 2632
rect 15148 2604 15512 2632
rect 15092 2576 15512 2604
rect 15848 2576 15988 2632
rect 17024 2604 17388 2632
rect 17920 2604 18480 2632
rect 17024 2576 17360 2604
rect 17920 2576 18368 2604
rect 15036 2548 15540 2576
rect 15820 2548 15988 2576
rect 17052 2548 17332 2576
rect 17920 2548 18256 2576
rect 14980 2520 15568 2548
rect 15792 2520 15960 2548
rect 17080 2520 17304 2548
rect 17920 2520 18144 2548
rect 14924 2492 15344 2520
rect 15400 2492 15624 2520
rect 15736 2492 15960 2520
rect 14868 2464 15288 2492
rect 15428 2464 15932 2492
rect 14812 2436 15232 2464
rect 15456 2436 15904 2464
rect 14756 2408 15176 2436
rect 15512 2408 15848 2436
rect 14700 2380 15120 2408
rect 15540 2380 15820 2408
rect 14644 2352 15064 2380
rect 14588 2324 15008 2352
rect 14532 2296 14952 2324
rect 14476 2268 14896 2296
rect 14420 2240 14840 2268
rect 14364 2212 14784 2240
rect 14308 2184 14728 2212
rect 14252 2156 14672 2184
rect 14196 2128 14616 2156
rect 14140 2100 14560 2128
rect 14084 2072 14504 2100
rect 14028 2044 14448 2072
rect 13972 2016 14392 2044
rect 13916 1988 14336 2016
rect 13860 1960 14280 1988
rect 13804 1932 14224 1960
rect 13748 1904 14168 1932
rect 13692 1876 14112 1904
rect 13636 1848 14056 1876
rect 13580 1820 14000 1848
rect 13524 1792 13944 1820
rect 13468 1764 13888 1792
rect 13384 1736 13832 1764
rect 13328 1708 13776 1736
rect 13272 1680 13720 1708
rect 13216 1652 13664 1680
rect 13160 1624 13608 1652
rect 13104 1596 13552 1624
rect 13048 1568 13496 1596
rect 7336 1540 7784 1568
rect 12768 1540 13440 1568
rect 1260 1512 1876 1540
rect 7112 1512 7728 1540
rect 12768 1512 13384 1540
rect 1260 1484 1820 1512
rect 7112 1484 7672 1512
rect 12768 1484 13328 1512
rect 1260 1456 1736 1484
rect 7112 1456 7616 1484
rect 12768 1456 13272 1484
rect 1260 1428 1680 1456
rect 7112 1428 7560 1456
rect 12768 1428 13216 1456
rect 1260 1400 1624 1428
rect 7112 1400 7504 1428
rect 12768 1400 13160 1428
rect 1260 1372 1568 1400
rect 7112 1372 7448 1400
rect 12768 1372 13104 1400
rect 1260 1344 1512 1372
rect 7112 1344 7392 1372
rect 12768 1344 13048 1372
rect 1260 1316 1456 1344
rect 7112 1316 7336 1344
rect 12768 1316 12992 1344
rect 1260 1288 1400 1316
rect 7112 1288 7280 1316
rect 12768 1288 12936 1316
rect 1260 1260 1344 1288
rect 7112 1260 7224 1288
rect 12768 1260 12880 1288
rect 1260 1232 1288 1260
rect 7112 1232 7168 1260
rect 12768 1232 12824 1260
rect 17136 140 17276 2520
rect 17920 2492 18032 2520
rect 0 0 17276 140
<< end >>
