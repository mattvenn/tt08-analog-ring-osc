magic
tech sky130A
magscale 1 2
timestamp 1725540246
<< error_p >>
rect -269 981 -211 987
rect -77 981 -19 987
rect 115 981 173 987
rect 307 981 365 987
rect -269 947 -257 981
rect -77 947 -65 981
rect 115 947 127 981
rect 307 947 319 981
rect -269 941 -211 947
rect -77 941 -19 947
rect 115 941 173 947
rect 307 941 365 947
rect -365 -947 -307 -941
rect -173 -947 -115 -941
rect 19 -947 77 -941
rect 211 -947 269 -941
rect -365 -981 -353 -947
rect -173 -981 -161 -947
rect 19 -981 31 -947
rect 211 -981 223 -947
rect -365 -987 -307 -981
rect -173 -987 -115 -981
rect 19 -987 77 -981
rect 211 -987 269 -981
<< nwell >>
rect -551 -1119 551 1119
<< pmos >>
rect -351 -900 -321 900
rect -255 -900 -225 900
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
rect 225 -900 255 900
rect 321 -900 351 900
<< pdiff >>
rect -413 888 -351 900
rect -413 -888 -401 888
rect -367 -888 -351 888
rect -413 -900 -351 -888
rect -321 888 -255 900
rect -321 -888 -305 888
rect -271 -888 -255 888
rect -321 -900 -255 -888
rect -225 888 -159 900
rect -225 -888 -209 888
rect -175 -888 -159 888
rect -225 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 225 900
rect 159 -888 175 888
rect 209 -888 225 888
rect 159 -900 225 -888
rect 255 888 321 900
rect 255 -888 271 888
rect 305 -888 321 888
rect 255 -900 321 -888
rect 351 888 413 900
rect 351 -888 367 888
rect 401 -888 413 888
rect 351 -900 413 -888
<< pdiffc >>
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
<< nsubdiff >>
rect -515 1049 -419 1083
rect 419 1049 515 1083
rect -515 987 -481 1049
rect 481 987 515 1049
rect -515 -1049 -481 -987
rect 481 -1049 515 -987
rect -515 -1083 -419 -1049
rect 419 -1083 515 -1049
<< nsubdiffcont >>
rect -419 1049 419 1083
rect -515 -987 -481 987
rect 481 -987 515 987
rect -419 -1083 419 -1049
<< poly >>
rect -273 981 -207 997
rect -273 947 -257 981
rect -223 947 -207 981
rect -273 931 -207 947
rect -81 981 -15 997
rect -81 947 -65 981
rect -31 947 -15 981
rect -81 931 -15 947
rect 111 981 177 997
rect 111 947 127 981
rect 161 947 177 981
rect 111 931 177 947
rect 303 981 369 997
rect 303 947 319 981
rect 353 947 369 981
rect 303 931 369 947
rect -351 900 -321 926
rect -255 900 -225 931
rect -159 900 -129 926
rect -63 900 -33 931
rect 33 900 63 926
rect 129 900 159 931
rect 225 900 255 926
rect 321 900 351 931
rect -351 -931 -321 -900
rect -255 -926 -225 -900
rect -159 -931 -129 -900
rect -63 -926 -33 -900
rect 33 -931 63 -900
rect 129 -926 159 -900
rect 225 -931 255 -900
rect 321 -926 351 -900
rect -369 -947 -303 -931
rect -369 -981 -353 -947
rect -319 -981 -303 -947
rect -369 -997 -303 -981
rect -177 -947 -111 -931
rect -177 -981 -161 -947
rect -127 -981 -111 -947
rect -177 -997 -111 -981
rect 15 -947 81 -931
rect 15 -981 31 -947
rect 65 -981 81 -947
rect 15 -997 81 -981
rect 207 -947 273 -931
rect 207 -981 223 -947
rect 257 -981 273 -947
rect 207 -997 273 -981
<< polycont >>
rect -257 947 -223 981
rect -65 947 -31 981
rect 127 947 161 981
rect 319 947 353 981
rect -353 -981 -319 -947
rect -161 -981 -127 -947
rect 31 -981 65 -947
rect 223 -981 257 -947
<< locali >>
rect -515 1049 -419 1083
rect 419 1049 515 1083
rect -515 987 -481 1049
rect 481 987 515 1049
rect -273 947 -257 981
rect -223 947 -207 981
rect -81 947 -65 981
rect -31 947 -15 981
rect 111 947 127 981
rect 161 947 177 981
rect 303 947 319 981
rect 353 947 369 981
rect -401 888 -367 904
rect -401 -904 -367 -888
rect -305 888 -271 904
rect -305 -904 -271 -888
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect 271 888 305 904
rect 271 -904 305 -888
rect 367 888 401 904
rect 367 -904 401 -888
rect -369 -981 -353 -947
rect -319 -981 -303 -947
rect -177 -981 -161 -947
rect -127 -981 -111 -947
rect 15 -981 31 -947
rect 65 -981 81 -947
rect 207 -981 223 -947
rect 257 -981 273 -947
rect -515 -1049 -481 -987
rect 481 -1049 515 -987
rect -515 -1083 -419 -1049
rect 419 -1083 515 -1049
<< viali >>
rect -257 947 -223 981
rect -65 947 -31 981
rect 127 947 161 981
rect 319 947 353 981
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect -353 -981 -319 -947
rect -161 -981 -127 -947
rect 31 -981 65 -947
rect 223 -981 257 -947
<< metal1 >>
rect -269 981 -211 987
rect -269 947 -257 981
rect -223 947 -211 981
rect -269 941 -211 947
rect -77 981 -19 987
rect -77 947 -65 981
rect -31 947 -19 981
rect -77 941 -19 947
rect 115 981 173 987
rect 115 947 127 981
rect 161 947 173 981
rect 115 941 173 947
rect 307 981 365 987
rect 307 947 319 981
rect 353 947 365 981
rect 307 941 365 947
rect -407 888 -361 900
rect -407 -888 -401 888
rect -367 -888 -361 888
rect -407 -900 -361 -888
rect -311 888 -265 900
rect -311 -888 -305 888
rect -271 -888 -265 888
rect -311 -900 -265 -888
rect -215 888 -169 900
rect -215 -888 -209 888
rect -175 -888 -169 888
rect -215 -900 -169 -888
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 169 888 215 900
rect 169 -888 175 888
rect 209 -888 215 888
rect 169 -900 215 -888
rect 265 888 311 900
rect 265 -888 271 888
rect 305 -888 311 888
rect 265 -900 311 -888
rect 361 888 407 900
rect 361 -888 367 888
rect 401 -888 407 888
rect 361 -900 407 -888
rect -365 -947 -307 -941
rect -365 -981 -353 -947
rect -319 -981 -307 -947
rect -365 -987 -307 -981
rect -173 -947 -115 -941
rect -173 -981 -161 -947
rect -127 -981 -115 -947
rect -173 -987 -115 -981
rect 19 -947 77 -941
rect 19 -981 31 -947
rect 65 -981 77 -947
rect 19 -987 77 -981
rect 211 -947 269 -941
rect 211 -981 223 -947
rect 257 -981 269 -947
rect 211 -987 269 -981
<< properties >>
string FIXED_BBOX -498 -1066 498 1066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9.0 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
