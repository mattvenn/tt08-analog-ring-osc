magic
tech sky130A
magscale 1 2
timestamp 1725540246
<< error_p >>
rect -269 372 -211 378
rect -77 372 -19 378
rect 115 372 173 378
rect 307 372 365 378
rect -269 338 -257 372
rect -77 338 -65 372
rect 115 338 127 372
rect 307 338 319 372
rect -269 332 -211 338
rect -77 332 -19 338
rect 115 332 173 338
rect 307 332 365 338
rect -365 -338 -307 -332
rect -173 -338 -115 -332
rect 19 -338 77 -332
rect 211 -338 269 -332
rect -365 -372 -353 -338
rect -173 -372 -161 -338
rect 19 -372 31 -338
rect 211 -372 223 -338
rect -365 -378 -307 -372
rect -173 -378 -115 -372
rect 19 -378 77 -372
rect 211 -378 269 -372
<< pwell >>
rect -551 -510 551 510
<< nmos >>
rect -351 -300 -321 300
rect -255 -300 -225 300
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
rect 225 -300 255 300
rect 321 -300 351 300
<< ndiff >>
rect -413 288 -351 300
rect -413 -288 -401 288
rect -367 -288 -351 288
rect -413 -300 -351 -288
rect -321 288 -255 300
rect -321 -288 -305 288
rect -271 -288 -255 288
rect -321 -300 -255 -288
rect -225 288 -159 300
rect -225 -288 -209 288
rect -175 -288 -159 288
rect -225 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 225 300
rect 159 -288 175 288
rect 209 -288 225 288
rect 159 -300 225 -288
rect 255 288 321 300
rect 255 -288 271 288
rect 305 -288 321 288
rect 255 -300 321 -288
rect 351 288 413 300
rect 351 -288 367 288
rect 401 -288 413 288
rect 351 -300 413 -288
<< ndiffc >>
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
<< psubdiff >>
rect -515 440 -419 474
rect 419 440 515 474
rect -515 378 -481 440
rect 481 378 515 440
rect -515 -440 -481 -378
rect 481 -440 515 -378
rect -515 -474 -419 -440
rect 419 -474 515 -440
<< psubdiffcont >>
rect -419 440 419 474
rect -515 -378 -481 378
rect 481 -378 515 378
rect -419 -474 419 -440
<< poly >>
rect -273 372 -207 388
rect -273 338 -257 372
rect -223 338 -207 372
rect -351 300 -321 326
rect -273 322 -207 338
rect -81 372 -15 388
rect -81 338 -65 372
rect -31 338 -15 372
rect -255 300 -225 322
rect -159 300 -129 326
rect -81 322 -15 338
rect 111 372 177 388
rect 111 338 127 372
rect 161 338 177 372
rect -63 300 -33 322
rect 33 300 63 326
rect 111 322 177 338
rect 303 372 369 388
rect 303 338 319 372
rect 353 338 369 372
rect 129 300 159 322
rect 225 300 255 326
rect 303 322 369 338
rect 321 300 351 322
rect -351 -322 -321 -300
rect -369 -338 -303 -322
rect -255 -326 -225 -300
rect -159 -322 -129 -300
rect -369 -372 -353 -338
rect -319 -372 -303 -338
rect -369 -388 -303 -372
rect -177 -338 -111 -322
rect -63 -326 -33 -300
rect 33 -322 63 -300
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect -177 -388 -111 -372
rect 15 -338 81 -322
rect 129 -326 159 -300
rect 225 -322 255 -300
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 15 -388 81 -372
rect 207 -338 273 -322
rect 321 -326 351 -300
rect 207 -372 223 -338
rect 257 -372 273 -338
rect 207 -388 273 -372
<< polycont >>
rect -257 338 -223 372
rect -65 338 -31 372
rect 127 338 161 372
rect 319 338 353 372
rect -353 -372 -319 -338
rect -161 -372 -127 -338
rect 31 -372 65 -338
rect 223 -372 257 -338
<< locali >>
rect -515 440 -419 474
rect 419 440 515 474
rect -515 378 -481 440
rect 481 378 515 440
rect -273 338 -257 372
rect -223 338 -207 372
rect -81 338 -65 372
rect -31 338 -15 372
rect 111 338 127 372
rect 161 338 177 372
rect 303 338 319 372
rect 353 338 369 372
rect -401 288 -367 304
rect -401 -304 -367 -288
rect -305 288 -271 304
rect -305 -304 -271 -288
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect 271 288 305 304
rect 271 -304 305 -288
rect 367 288 401 304
rect 367 -304 401 -288
rect -369 -372 -353 -338
rect -319 -372 -303 -338
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 207 -372 223 -338
rect 257 -372 273 -338
rect -515 -440 -481 -378
rect 481 -440 515 -378
rect -515 -474 -419 -440
rect 419 -474 515 -440
<< viali >>
rect -257 338 -223 372
rect -65 338 -31 372
rect 127 338 161 372
rect 319 338 353 372
rect -401 -288 -367 288
rect -305 -288 -271 288
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect 271 -288 305 288
rect 367 -288 401 288
rect -353 -372 -319 -338
rect -161 -372 -127 -338
rect 31 -372 65 -338
rect 223 -372 257 -338
<< metal1 >>
rect -269 372 -211 378
rect -269 338 -257 372
rect -223 338 -211 372
rect -269 332 -211 338
rect -77 372 -19 378
rect -77 338 -65 372
rect -31 338 -19 372
rect -77 332 -19 338
rect 115 372 173 378
rect 115 338 127 372
rect 161 338 173 372
rect 115 332 173 338
rect 307 372 365 378
rect 307 338 319 372
rect 353 338 365 372
rect 307 332 365 338
rect -407 288 -361 300
rect -407 -288 -401 288
rect -367 -288 -361 288
rect -407 -300 -361 -288
rect -311 288 -265 300
rect -311 -288 -305 288
rect -271 -288 -265 288
rect -311 -300 -265 -288
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect 265 288 311 300
rect 265 -288 271 288
rect 305 -288 311 288
rect 265 -300 311 -288
rect 361 288 407 300
rect 361 -288 367 288
rect 401 -288 407 288
rect 361 -300 407 -288
rect -365 -338 -307 -332
rect -365 -372 -353 -338
rect -319 -372 -307 -338
rect -365 -378 -307 -372
rect -173 -338 -115 -332
rect -173 -372 -161 -338
rect -127 -372 -115 -338
rect -173 -378 -115 -372
rect 19 -338 77 -332
rect 19 -372 31 -338
rect 65 -372 77 -338
rect 19 -378 77 -372
rect 211 -338 269 -332
rect 211 -372 223 -338
rect 257 -372 269 -338
rect 211 -378 269 -372
<< properties >>
string FIXED_BBOX -498 -457 498 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
