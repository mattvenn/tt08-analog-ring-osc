MACRO tt_um_mattvenn_analog_ring_osc
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_analog_ring_osc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.000 BY 1.000 ;
END tt_um_mattvenn_analog_ring_osc
END LIBRARY

