magic
tech sky130A
magscale 1 2
timestamp 1725561929
<< nwell >>
rect 2640 136 3410 360
rect 2980 100 3410 136
rect 2980 40 3000 100
<< viali >>
rect 630 -10 664 24
rect 810 0 844 34
rect 906 -10 940 24
rect 1086 0 1120 34
rect 1182 -10 1216 24
rect 1362 0 1396 34
rect 1458 -10 1492 24
rect 1638 0 1672 34
rect 1734 -10 1768 24
rect 1914 0 1948 34
rect 2010 -10 2044 24
rect 2190 0 2224 34
rect 2286 -10 2320 24
rect 2466 0 2500 34
rect 2562 -10 2596 24
rect 2742 0 2776 34
rect 2830 -10 2864 24
rect 710 -484 744 -450
rect 890 -474 924 -440
rect 986 -484 1020 -450
rect 1166 -474 1200 -440
rect 1262 -484 1296 -450
rect 1442 -474 1476 -440
rect 1538 -484 1572 -450
rect 1718 -474 1752 -440
rect 1814 -484 1848 -450
rect 1994 -474 2028 -440
rect 2090 -484 2124 -450
rect 2270 -474 2304 -440
rect 2366 -484 2400 -450
rect 2546 -474 2580 -440
rect 2642 -484 2676 -450
rect 2822 -474 2856 -440
rect 2918 -484 2952 -450
<< metal1 >>
rect -200 600 3980 640
rect -200 420 260 600
rect 3020 420 3980 600
rect 4360 495 4640 640
rect -200 280 3980 420
rect 4240 425 4640 495
rect 4240 230 4310 425
rect 4360 280 4640 425
rect 3660 160 4310 230
rect 3660 120 3730 160
rect 3890 60 4440 70
rect -26 -10 -20 50
rect 40 -10 92 50
rect 620 34 860 50
rect 620 24 810 34
rect 620 -10 630 24
rect 664 0 810 24
rect 844 0 860 34
rect 664 -10 860 0
rect 620 -30 860 -10
rect 896 34 1136 50
rect 896 24 1086 34
rect 896 -10 906 24
rect 940 0 1086 24
rect 1120 0 1136 34
rect 940 -10 1136 0
rect 896 -30 1136 -10
rect 1172 34 1412 50
rect 1172 24 1362 34
rect 1172 -10 1182 24
rect 1216 0 1362 24
rect 1396 0 1412 34
rect 1216 -10 1412 0
rect 1172 -30 1412 -10
rect 1448 34 1688 50
rect 1448 24 1638 34
rect 1448 -10 1458 24
rect 1492 0 1638 24
rect 1672 0 1688 34
rect 1492 -10 1688 0
rect 1448 -30 1688 -10
rect 1724 34 1964 50
rect 1724 24 1914 34
rect 1724 -10 1734 24
rect 1768 0 1914 24
rect 1948 0 1964 34
rect 1768 -10 1964 0
rect 1724 -30 1964 -10
rect 2000 34 2240 50
rect 2000 24 2190 34
rect 2000 -10 2010 24
rect 2044 0 2190 24
rect 2224 0 2240 34
rect 2044 -10 2240 0
rect 2000 -30 2240 -10
rect 2276 34 2516 50
rect 2276 24 2466 34
rect 2276 -10 2286 24
rect 2320 0 2466 24
rect 2500 0 2516 34
rect 2320 -10 2516 0
rect 2276 -30 2516 -10
rect 2552 34 2792 50
rect 2552 24 2742 34
rect 2552 -10 2562 24
rect 2596 0 2742 24
rect 2776 0 2792 34
rect 2596 -10 2792 0
rect 2552 -30 2792 -10
rect 2820 24 3060 50
rect 2820 -10 2830 24
rect 2864 -10 3060 24
rect 3840 0 3900 60
rect 3960 0 4440 60
rect 3890 -10 4440 0
rect 2820 -30 3060 -10
rect 4280 -160 4440 -10
rect -220 -204 276 -160
rect -220 -272 3980 -204
rect -220 -440 276 -272
rect 694 -440 934 -420
rect 694 -450 890 -440
rect 694 -484 710 -450
rect 744 -474 890 -450
rect 924 -474 934 -440
rect 744 -484 934 -474
rect 694 -500 934 -484
rect 970 -440 1210 -420
rect 970 -450 1166 -440
rect 970 -484 986 -450
rect 1020 -474 1166 -450
rect 1200 -474 1210 -440
rect 1020 -484 1210 -474
rect 970 -500 1210 -484
rect 1246 -440 1486 -420
rect 1246 -450 1442 -440
rect 1246 -484 1262 -450
rect 1296 -474 1442 -450
rect 1476 -474 1486 -440
rect 1296 -484 1486 -474
rect 1246 -500 1486 -484
rect 1522 -440 1762 -420
rect 1522 -450 1718 -440
rect 1522 -484 1538 -450
rect 1572 -474 1718 -450
rect 1752 -474 1762 -440
rect 1572 -484 1762 -474
rect 1522 -500 1762 -484
rect 1798 -440 2038 -420
rect 1798 -450 1994 -440
rect 1798 -484 1814 -450
rect 1848 -474 1994 -450
rect 2028 -474 2038 -440
rect 1848 -484 2038 -474
rect 1798 -500 2038 -484
rect 2074 -440 2314 -420
rect 2074 -450 2270 -440
rect 2074 -484 2090 -450
rect 2124 -474 2270 -450
rect 2304 -474 2314 -440
rect 2124 -484 2314 -474
rect 2074 -500 2314 -484
rect 2350 -440 2590 -420
rect 2350 -450 2546 -440
rect 2350 -484 2366 -450
rect 2400 -474 2546 -450
rect 2580 -474 2590 -440
rect 2400 -484 2590 -474
rect 2350 -500 2590 -484
rect 2626 -440 2866 -420
rect 2626 -450 2822 -440
rect 2626 -484 2642 -450
rect 2676 -474 2822 -450
rect 2856 -474 2866 -440
rect 2676 -484 2866 -474
rect 2626 -500 2866 -484
rect 2902 -450 3128 -420
rect 4280 -440 4640 -160
rect 2902 -484 2918 -450
rect 2952 -484 3128 -450
rect 2902 -500 3128 -484
rect -26 -650 -20 -590
rect 40 -600 170 -590
rect 40 -650 184 -600
rect 3340 -680 3900 -620
rect 3960 -680 3966 -620
rect -184 -880 3956 -748
rect -200 -1020 3980 -880
rect -200 -1200 260 -1020
rect 3020 -1200 3980 -1020
rect -200 -1240 3980 -1200
<< via1 >>
rect 260 420 3020 600
rect -20 -10 40 50
rect 3900 0 3960 60
rect -20 -650 40 -590
rect 3900 -680 3960 -620
rect 260 -1200 3020 -1020
<< metal2 >>
rect 200 600 3080 640
rect 200 420 260 600
rect 3020 420 3080 600
rect -20 50 40 56
rect -20 -590 40 -10
rect -20 -656 40 -650
rect 200 -880 3080 420
rect 3890 60 3970 70
rect 3890 0 3900 60
rect 3960 0 3970 60
rect 3890 -10 3970 0
rect 3900 -620 3960 -10
rect 3900 -686 3960 -680
rect -200 -1020 3080 -880
rect -200 -1200 260 -1020
rect 3020 -1200 3080 -1020
rect -200 -1240 3080 -1200
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1704896540
transform 1 0 2430 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1704896540
transform 1 0 498 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1704896540
transform 1 0 774 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1704896540
transform 1 0 1050 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1704896540
transform 1 0 1326 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1704896540
transform 1 0 1602 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1704896540
transform 1 0 1878 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1704896540
transform 1 0 2154 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1704896540
transform -1 0 774 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_9
timestamp 1704896540
transform 1 0 2706 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_10
timestamp 1704896540
transform -1 0 2982 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_11
timestamp 1704896540
transform -1 0 2706 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_12
timestamp 1704896540
transform -1 0 2430 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_13
timestamp 1704896540
transform -1 0 2154 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_14
timestamp 1704896540
transform -1 0 1878 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_15
timestamp 1704896540
transform -1 0 1602 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_16
timestamp 1704896540
transform -1 0 1326 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_17
timestamp 1704896540
transform -1 0 1050 0 -1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_0
timestamp 1704896540
transform 1 0 3350 0 1 -224
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1704896540
transform 1 0 18 0 -1 -388
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1704896540
transform 1 0 18 0 1 -212
box -38 -48 130 592
<< labels >>
flabel metal1 -220 -440 -20 -160 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 -200 280 -40 640 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal1 4360 280 4640 640 0 FreeSans 1600 0 0 0 enable
port 3 nsew
flabel metal1 4360 -440 4640 -160 0 FreeSans 1600 0 0 0 out
port 5 nsew
<< end >>
