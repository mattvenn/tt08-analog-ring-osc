magic
tech sky130A
magscale 1 2
timestamp 1725561279
<< nwell >>
rect 2640 136 3410 360
rect 2980 100 3410 136
rect 2980 40 3000 100
<< viali >>
rect 630 -10 664 24
rect 810 0 844 34
rect 906 -10 940 24
rect 1086 0 1120 34
rect 1182 -10 1216 24
rect 1362 0 1396 34
rect 1458 -10 1492 24
rect 1638 0 1672 34
rect 1734 -10 1768 24
rect 1914 0 1948 34
rect 2010 -10 2044 24
rect 2190 0 2224 34
rect 2286 -10 2320 24
rect 2466 0 2500 34
rect 2562 -10 2596 24
rect 2742 0 2776 34
rect 2830 -10 2864 24
rect 710 -620 744 -586
rect 890 -610 924 -576
rect 986 -620 1020 -586
rect 1166 -610 1200 -576
rect 1262 -620 1296 -586
rect 1442 -610 1476 -576
rect 1538 -620 1572 -586
rect 1718 -610 1752 -576
rect 1814 -620 1848 -586
rect 1994 -610 2028 -576
rect 2090 -620 2124 -586
rect 2270 -610 2304 -576
rect 2366 -620 2400 -586
rect 2546 -610 2580 -576
rect 2642 -620 2676 -586
rect 2822 -610 2856 -576
rect 2918 -620 2952 -586
<< metal1 >>
rect -200 600 3980 640
rect -200 420 260 600
rect 3020 420 3980 600
rect 4360 495 4640 640
rect -200 280 3980 420
rect 4240 425 4640 495
rect 4240 230 4310 425
rect 4360 280 4640 425
rect 3660 160 4310 230
rect 3660 120 3730 160
rect 3890 60 4440 70
rect -26 -10 -20 50
rect 40 -10 92 50
rect 620 34 860 50
rect 620 24 810 34
rect 620 -10 630 24
rect 664 0 810 24
rect 844 0 860 34
rect 664 -10 860 0
rect 620 -30 860 -10
rect 896 34 1136 50
rect 896 24 1086 34
rect 896 -10 906 24
rect 940 0 1086 24
rect 1120 0 1136 34
rect 940 -10 1136 0
rect 896 -30 1136 -10
rect 1172 34 1412 50
rect 1172 24 1362 34
rect 1172 -10 1182 24
rect 1216 0 1362 24
rect 1396 0 1412 34
rect 1216 -10 1412 0
rect 1172 -30 1412 -10
rect 1448 34 1688 50
rect 1448 24 1638 34
rect 1448 -10 1458 24
rect 1492 0 1638 24
rect 1672 0 1688 34
rect 1492 -10 1688 0
rect 1448 -30 1688 -10
rect 1724 34 1964 50
rect 1724 24 1914 34
rect 1724 -10 1734 24
rect 1768 0 1914 24
rect 1948 0 1964 34
rect 1768 -10 1964 0
rect 1724 -30 1964 -10
rect 2000 34 2240 50
rect 2000 24 2190 34
rect 2000 -10 2010 24
rect 2044 0 2190 24
rect 2224 0 2240 34
rect 2044 -10 2240 0
rect 2000 -30 2240 -10
rect 2276 34 2516 50
rect 2276 24 2466 34
rect 2276 -10 2286 24
rect 2320 0 2466 24
rect 2500 0 2516 34
rect 2320 -10 2516 0
rect 2276 -30 2516 -10
rect 2552 34 2792 50
rect 2552 24 2742 34
rect 2552 -10 2562 24
rect 2596 0 2742 24
rect 2776 0 2792 34
rect 2596 -10 2792 0
rect 2552 -30 2792 -10
rect 2820 24 3060 50
rect 2820 -10 2830 24
rect 2864 -10 3060 24
rect 3840 0 3900 60
rect 3960 0 4440 60
rect 3890 -10 4440 0
rect 2820 -30 3060 -10
rect 4280 -160 4440 -10
rect -220 -440 3980 -160
rect 4280 -440 4640 -160
rect 694 -576 934 -556
rect 694 -586 890 -576
rect -26 -650 -20 -590
rect 40 -600 170 -590
rect 40 -650 184 -600
rect 694 -620 710 -586
rect 744 -610 890 -586
rect 924 -610 934 -576
rect 744 -620 934 -610
rect 694 -636 934 -620
rect 970 -576 1210 -556
rect 970 -586 1166 -576
rect 970 -620 986 -586
rect 1020 -610 1166 -586
rect 1200 -610 1210 -576
rect 1020 -620 1210 -610
rect 970 -636 1210 -620
rect 1246 -576 1486 -556
rect 1246 -586 1442 -576
rect 1246 -620 1262 -586
rect 1296 -610 1442 -586
rect 1476 -610 1486 -576
rect 1296 -620 1486 -610
rect 1246 -636 1486 -620
rect 1522 -576 1762 -556
rect 1522 -586 1718 -576
rect 1522 -620 1538 -586
rect 1572 -610 1718 -586
rect 1752 -610 1762 -576
rect 1572 -620 1762 -610
rect 1522 -636 1762 -620
rect 1798 -576 2038 -556
rect 1798 -586 1994 -576
rect 1798 -620 1814 -586
rect 1848 -610 1994 -586
rect 2028 -610 2038 -576
rect 1848 -620 2038 -610
rect 1798 -636 2038 -620
rect 2074 -576 2314 -556
rect 2074 -586 2270 -576
rect 2074 -620 2090 -586
rect 2124 -610 2270 -586
rect 2304 -610 2314 -576
rect 2124 -620 2314 -610
rect 2074 -636 2314 -620
rect 2350 -576 2590 -556
rect 2350 -586 2546 -576
rect 2350 -620 2366 -586
rect 2400 -610 2546 -586
rect 2580 -610 2590 -576
rect 2400 -620 2590 -610
rect 2350 -636 2590 -620
rect 2626 -576 2866 -556
rect 2626 -586 2822 -576
rect 2626 -620 2642 -586
rect 2676 -610 2822 -586
rect 2856 -610 2866 -576
rect 2676 -620 2866 -610
rect 2626 -636 2866 -620
rect 2902 -586 3142 -556
rect 2902 -620 2918 -586
rect 2952 -620 3142 -586
rect 2902 -636 3142 -620
rect 3340 -680 3900 -620
rect 3960 -680 3966 -620
rect -200 -1020 3980 -880
rect -200 -1200 260 -1020
rect 3020 -1200 3980 -1020
rect -200 -1240 3980 -1200
<< via1 >>
rect 260 420 3020 600
rect -20 -10 40 50
rect 3900 0 3960 60
rect -20 -650 40 -590
rect 3900 -680 3960 -620
rect 260 -1200 3020 -1020
<< metal2 >>
rect 200 600 3080 640
rect 200 420 260 600
rect 3020 420 3080 600
rect -20 50 40 56
rect -20 -590 40 -10
rect -20 -656 40 -650
rect 200 -880 3080 420
rect 3890 60 3970 70
rect 3890 0 3900 60
rect 3960 0 3970 60
rect 3890 -10 3970 0
rect 3900 -620 3960 -10
rect 3900 -686 3960 -680
rect -200 -1020 3080 -880
rect -200 -1200 260 -1020
rect 3020 -1200 3080 -1020
rect -200 -1240 3080 -1200
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1704896540
transform 1 0 2430 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1704896540
transform 1 0 498 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1704896540
transform 1 0 774 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1704896540
transform 1 0 1050 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1704896540
transform 1 0 1326 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1704896540
transform 1 0 1602 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1704896540
transform 1 0 1878 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1704896540
transform 1 0 2154 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1704896540
transform -1 0 774 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_9
timestamp 1704896540
transform 1 0 2706 0 1 -224
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_10
timestamp 1704896540
transform -1 0 2982 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_11
timestamp 1704896540
transform -1 0 2706 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_12
timestamp 1704896540
transform -1 0 2430 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_13
timestamp 1704896540
transform -1 0 2154 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_14
timestamp 1704896540
transform -1 0 1878 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_15
timestamp 1704896540
transform -1 0 1602 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_16
timestamp 1704896540
transform -1 0 1326 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_17
timestamp 1704896540
transform -1 0 1050 0 -1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  sky130_fd_sc_hd__nand2_2_0
timestamp 1704896540
transform 1 0 3350 0 1 -224
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1704896540
transform 1 0 18 0 -1 -388
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1704896540
transform 1 0 18 0 1 -212
box -38 -48 130 592
<< labels >>
flabel metal1 -220 -440 -20 -160 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 -200 280 -40 640 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal1 4360 280 4640 640 0 FreeSans 1600 0 0 0 enable
port 3 nsew
flabel metal1 4360 -440 4640 -160 0 FreeSans 1600 0 0 0 out
port 5 nsew
<< end >>
